`ifndef   _fifo_vh_
  `define _fifo_vh_

  `define DATA_WIDTH 32
  
`endif